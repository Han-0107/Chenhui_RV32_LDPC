
`timescale 1 ns/ 1 ps
module ldpc_encoder(
	clk,
	rst_n,
	msg,
	code,
	tx_en,
	uart_done
	);

	input  		  clk;													// ????? 50MHz
	input  		  rst_n;												// ??λ??????????Ч
	input  		  uart_done;
	output         tx_en;
	input  [3:0]  msg;													// ??????? 
	output [11:0] code;													// ???????? 
reg [3:0]     msg_r;
    /*********************************************************************************************
    //  ????????LDPC???????
    //  ??????????????????н???LDPC????
	//			   ????(8??12)???????????LDPC???????0.33???????3??4???????2??3 	 
    //             ????????????????????????У??????c??????????????????code            
	//   			| 0	 0	1	0	0	1	0	0	1	0	1	0 |
	//				| 0	 1	0	0	0	1	0	0	0	0	0	1 |
	//  			| 0	 1	0	0	0	0	1	0	0	0	1	0 |
	//  У?????H=  | 0	 0	0	1	1	1	0	0	0	1	0	0 |       ??code*H'=0 ??code??? ????????msg
	//  			| 0	 0	0	1	0	0	0	1	1	0	0	1 |
	//  			| 1	 0	0	0	1	0	0	0	0	0	0	0 |
	//  			| 1	 0	1	0	0	0	1	1	0	0	0	0 |
	//   			| 0	 1	1	0	0	0	0	0	0	1	0	0 |
	//		 	                 
	//                          ??????
    //  ??H=[A | B] ???? [I | P] ??I???λ???? 
    //  ??u????????? u=[c | s]  s???????? c?У??????
    //  ???  H*u' = u*H' = 0
    //  ??????
	//			 _    _
	//			 | c' |
	//	  [I | P]|    | = 0
	//			 | s' |
	//			 -    -
	//	 I*c' + P*s' = 0
	//	 I*c' = P*s' (??GF(2)??) ->  I*c'=-P*s' 
	//   ?????GF(2)???? P*s'+ P*s'=0 ???? P*s'=-P*s' I*c' = P*s' ->   c'=I'*P*s' =P*s' -> c' = P*s' 
	//	 ????u=[c | s]?????????????????
	//	 ??????????????н??????н?????
	//	 ????????н???col_recoeder??????????????????????????????н??????ɡ?
	//	 ??????????u????????н??????u=[c | s]?????沿??s??????????????????С?
	//   
	//   ????У?????H?????????????????H??????[I | P]??P?8??6?е?????????P??????н???col_recoeder????????
	//     | 1 1 1 0 |
	//	p= | 0 1 0 1 |      col_recoeder= |0 0 0 0 0 0 0 9| ??0????任??
	//     | 0 0 0 1 |
	//     | 1 1 1 0 |
	//	   | 1 1 1 0 |
	//     | 0 1 0 0 |
	//     | 0 1 1 1 |
	//     | 0 1 1 1 |
    //*********************************************************************************************/	

always@(posedge clk or negedge rst_n)
	begin
	   if(!rst_n)
	       msg_r <= 0;
	   else if(uart_done)
	       msg_r <= msg;
	   else
	      msg_r <= msg_r;
	end

	// ?????? ???????????У????????? ???????? ?????б任??? ????????????
	reg [1:0] clk_count;
	reg        tx_flag;
	
	always@(posedge clk or negedge rst_n)
	   if(!rst_n)
	       tx_flag <= 0;
	   else if(uart_done)
	       tx_flag <= 1;
	   else if(clk_count==2'd3)
	       tx_flag <= 0;
	   else
	       tx_flag <= tx_flag;
	  
	always@(posedge clk or negedge rst_n)
	begin
		if(rst_n == 2'b00)												//??λ?????Ч
			clk_count <= #1 2'b00;
		else if(tx_flag)
			clk_count <= #1 clk_count + 1'b1;
	   else
	       clk_count <= 2'd0;
	end
	
	
	// msg_r??P??????????? ???У??????
	reg [7:0] check;													// У??????
	always@(posedge clk or negedge rst_n)
	begin
		if(rst_n == 1'b0)
			check     <= #1 8'b0;
		else
		begin
			if(clk_count == 2'd1)
			begin														// msg??P??????????? ???У??????								
				check[7]  <= #1 msg_r[3]+msg_r[2]+msg_r[1];
				check[6]  <= #1 msg_r[2]+msg_r[0];
				check[5]  <= #1 msg_r[0];
				check[4]  <= #1 msg_r[3]+msg_r[2]+msg_r[1];
				check[3]  <= #1 msg_r[3]+msg_r[2]+msg_r[1];
				check[2]  <= #1 msg_r[2];
				check[1]  <= #1 msg_r[2]+msg_r[1]+msg_r[0];
				check[0]  <= #1 msg_r[2]+msg_r[1]+msg_r[0];
			end
			else
				check <= #1 8'b0;
		end
	end
	
	// ?????б任?????????????????	|0 0 0 0 0 0 0 9|  u=[c | s] 
	reg [11:0] code;													
	always@(posedge clk or negedge rst_n)
	begin
		if(rst_n == 1'b0)
			code <= #1 12'b0;
			
		else
		begin
			if(clk_count == 2'd2)
				code <= #1 {check[7:1],msg_r[3],check[0],msg_r[2:0]}; 	// ???е?8λ???9λ???н??? ????????? ???????????????	
																	// ??????????????????????е?8??9λ????	
			else
				code  <= #1 code;			
		end
	end	
	
	assign     tx_en = (clk_count == 2'd3)?1'b1:1'b0;
	
endmodule

//LDPC????????????
//?????H???????????LDPC??????????H???????????????LDPC?????????
//?????H??????б任?????[I | P]?????У?I?8*8???λ????P?4*8?????
//???????????????????P?????У?????c???????s????
//			 _    _
//			 | c' |
//	  [I | P]|    | = 0
//			 | s' |
//			 -    -
//????????????c??s????????P???????γ?????У???????????б任????????????????????code???????????????任??????????????????H????????????????????б任??????
//??????code